library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity test_memory_only is
end test_memory_only;

architecture tb of test_memory_only is
    
    signal clk : std_logic := '0';
    signal write_enable : std_logic := '0';
    signal read_enable : std_logic := '0';
    signal address : unsigned(11 downto 0) := (others => '0');
    signal bus_input : std_logic_vector(15 downto 0) := (others => '0');
    signal bus_output : std_logic_vector(15 downto 0);
    
begin
    
    clk <= not clk after 10 ns;
    
    MEM: entity work.memory
    port map(
        clk => clk,
        write_enable => write_enable,
        read_enable => read_enable,
        address => address,
        bus_input => bus_input,
        bus_output => bus_output
    );
    
    process
    begin
        
        report "??? ?????";
        wait for 20 ns;
        
        address <= "000000000000";
        bus_input <= "0000010000010100";
        write_enable <= '1';
        wait for 20 ns;
        write_enable <= '0';
        wait for 20 ns;
        
        report "????? ?? ???? 0";
        
        read_enable <= '1';
        wait for 20 ns;
        
        if bus_output = "0000010000010100" then
            report "?????? ????";
        else
            report "?????? ??????";
        end if;
        
        read_enable <= '0';
        wait for 20 ns;
        
        address <= "000000000001";
        bus_input <= "0000000000001111";
        write_enable <= '1';
        wait for 20 ns;
        write_enable <= '0';
        wait for 20 ns;
        
        address <= "000000000001";
        read_enable <= '1';
        wait for 20 ns;
        
        if bus_output = "0000000000001111" then
            report "?????? ?? ???? 1 ????";
        else
            report "?????? ?? ???? 1 ??????";
        end if;
        
        read_enable <= '0';
        wait for 20 ns;
        
        address <= "000000000000";
        read_enable <= '1';
        wait for 20 ns;
        
        if bus_output = "0000010000010100" then
            report "???????? ????";
        else
            report "???????? ??????";
        end if;
        
        read_enable <= '0';
        
        report "????? ???";
        wait;
        
    end process;
    
end tb;
